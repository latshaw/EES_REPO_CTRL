LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TEMP_LIMIT_COEFF IS

	PORT(JMPR_SET : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 TEMP_LIMIT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
		 );
		 
END ENTITY TEMP_LIMIT_COEFF;

ARCHITECTURE BEHAVIOR OF TEMP_LIMIT_COEFF IS

BEGIN


TEMP_LIMIT <= x"01FF" WHEN JMPR_SET = "000" ELSE
			  x"03FF" WHEN JMPR_SET = "001" ELSE
			  x"05FF" WHEN JMPR_SET = "010" ELSE
			  x"07FF" WHEN JMPR_SET = "011" ELSE
			  x"09FF" WHEN JMPR_SET = "100" ELSE
			  x"0BFF" WHEN JMPR_SET = "101" ELSE
			  x"0DFF" WHEN JMPR_SET = "110" ELSE
			  x"0FFF";


END ARCHITECTURE BEHAVIOR;