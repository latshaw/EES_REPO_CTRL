LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE WORK.COMPONENTS.ALL;

ENTITY MCP3202 IS
	PORT(CLOCK : IN STD_LOGIC;
		 RESET : IN STD_LOGIC;
		 HTR_ADC_DO : IN STD_LOGIC;
		 
		 HTR_CURRENT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 HTR_VOLTAGE : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 HTR_ADC_CLK : OUT STD_LOGIC;
		 HTR_ADC_DI : OUT STD_LOGIC;
		 HTR_ADC_CS : OUT STD_LOGIC
		 
		 
		 );
END ENTITY MCP3202;

ARCHITECTURE BEHAVIOR OF MCP3202 IS

SIGNAL EN_ADC_DATA			: STD_LOGIC;
SIGNAL ADC_DATA				: STD_LOGIC_VECTOR(11 DOWNTO 0);

SIGNAL EN_ADC_CNTRL			: STD_LOGIC;
SIGNAL LD_ADC_CNTRL			: STD_LOGIC;
SIGNAL INP_ADC_CNTRL		: STD_LOGIC_VECTOR(15 DOWNTO 0);

SIGNAL CLR_BIT_COUNT		: STD_LOGIC;
SIGNAL EN_BIT_COUNT			: STD_LOGIC;
SIGNAL BIT_COUNT			: STD_LOGIC_VECTOR(4 DOWNTO 0);

SIGNAL CLR_CLK_COUNT		: STD_LOGIC;
SIGNAL EN_CLK_COUNT			: STD_LOGIC;
SIGNAL CLK_COUNT			: STD_LOGIC_VECTOR(5 DOWNTO 0);

SIGNAL EN_CHNL_COUNT		: STD_LOGIC;
SIGNAL CHNL_COUNT			: STD_LOGIC_VECTOR(1 DOWNTO 0);

SIGNAL EN_HTRI				: STD_LOGIC;
SIGNAL HTR_I_TEMP			: STD_LOGIC_VECTOR(11 DOWNTO 0);

SIGNAL EN_HTRV				: STD_LOGIC;
SIGNAL HTR_V_TEMP			: STD_LOGIC_VECTOR(11 DOWNTO 0);


SIGNAL ONE					: STD_LOGIC;

TYPE STATE_TYPE IS (INIT, CS_HIGH, CS_LOW, CLK_LOW, CLK_HIGH, DONE);
SIGNAL STATE				: STATE_TYPE;



BEGIN

	ONE <= '1';
	
	
	HTR_I_REG: REGNE
		GENERIC MAP(N => 12)
		PORT MAP(CLOCK	=> CLOCK, 
				 RESET	=> RESET,
				 CLEAR 	=> ONE,
				 EN		=> EN_HTRI,
				 INPUT	=> ADC_DATA,
				 OUTPUT	=> HTR_I_TEMP
				);	
				
	HTR_CURRENT <= "0000" & HTR_I_TEMP;
	EN_HTRI <= '1' WHEN STATE = DONE AND CHNL_COUNT (0) = '1' ELSE '0';
	
	HTR_V_REG: REGNE
		GENERIC MAP(N => 12)
		PORT MAP(CLOCK	=> CLOCK, 
				 RESET	=> RESET,
				 CLEAR 	=> ONE,
				 EN		=> EN_HTRV,
				 INPUT	=> ADC_DATA,
				 OUTPUT	=> HTR_V_TEMP
				);
				
	HTR_VOLTAGE <= "0000" & HTR_V_TEMP;
	EN_HTRV <= '1' WHEN STATE = DONE AND CHNL_COUNT (0) = '0' ELSE '0';
		

	ADC_CONV_DATA: SHIFT_LEFT_REG
		GENERIC MAP(N => 12)
		PORT MAP(CLOCK	=> CLOCK,
				 RESET	=> RESET,
				 EN		=> EN_ADC_DATA,
				 INP	=> HTR_ADC_DO,
				 OUTPUT	=> ADC_DATA
				);

	ADC_CNTRL_DATA: SHIFT_REG
		GENERIC MAP(N => 16)
		PORT MAP(CLOCK	=> CLOCK,
				 RESET	=> RESET,
				 EN		=> EN_ADC_CNTRL,
				 LOAD	=> LD_ADC_CNTRL,
				 INP	=> INP_ADC_CNTRL,
				 OUTPUT	=> HTR_ADC_DI
				);
				
	INP_ADC_CNTRL <= x"E000" WHEN CHNL_COUNT(0) = '1' ELSE x"C000";


	BIT_COUNTER: COUNTER
		GENERIC MAP(N => 5)
		PORT MAP(CLOCK	=> CLOCK,
				 RESET	=> RESET,
				 CLEAR	=> CLR_BIT_COUNT,
				 ENABLE	=> EN_BIT_COUNT,
				 COUNT	=> BIT_COUNT
				);

	CHNL_COUNTER: COUNTER
		GENERIC MAP(N => 2)
		PORT MAP(CLOCK	=> CLOCK,
				 RESET	=> RESET,
				 CLEAR	=> ONE,
				 ENABLE	=> EN_CHNL_COUNT,
				 COUNT	=> CHNL_COUNT
				);				

	CLOCK_COUNTER: COUNTER
		GENERIC MAP(N => 6)
		PORT MAP(CLOCK	=> CLOCK,
				 RESET	=> RESET,
				 CLEAR	=> CLR_CLK_COUNT,
				 ENABLE	=> EN_CLK_COUNT,
				 COUNT	=> CLK_COUNT
				);
				
				
				
	PROCESS(CLOCK, RESET)
	BEGIN
	
		IF(RESET = '0') THEN
			STATE <= INIT;
		ELSIF(CLOCK = '1' AND CLOCK'EVENT) THEN
			
			CASE STATE IS
			
				WHEN INIT => STATE <= CS_HIGH;
				
				WHEN CS_HIGH => IF CLK_COUNT = "110010" THEN STATE <= CS_LOW;
								ELSE STATE <= CS_HIGH;
								END IF;
								
				WHEN CS_LOW => STATE <= CLK_LOW;
				
				WHEN CLK_LOW => IF CLK_COUNT = "011000" THEN STATE <= CLK_HIGH;
								ELSE STATE <= CLK_LOW;
								END IF;
								
				WHEN CLK_HIGH => IF CLK_COUNT = "110001" THEN
									IF BIT_COUNT = "10000" THEN STATE <= DONE;
									ELSE STATE <= CLK_LOW;
									END IF;
								 ELSE STATE <= CLK_HIGH;
								 END IF;
								 
				WHEN DONE => STATE <= CS_HIGH;
				
			END CASE;
		END IF;
	END PROCESS;
						

	LD_ADC_CNTRL <= '1' WHEN STATE = INIT OR STATE = DONE ELSE '0';
	EN_ADC_CNTRL <= '1' WHEN (STATE = CLK_LOW AND CLK_COUNT = "000011" AND BIT_COUNT /= "00000") ELSE '0';
	
	EN_ADC_DATA <= '1' WHEN STATE = CLK_HIGH AND CLK_COUNT = "011011" ELSE '0'; 
	
	EN_CHNL_COUNT <= '1' WHEN (STATE = DONE) ELSE '0';

	EN_BIT_COUNT <= '1' WHEN STATE = CLK_HIGH AND CLK_COUNT = "110001" AND BIT_COUNT /= "10000" ELSE '0';
	CLR_BIT_COUNT <= '0' WHEN STATE = DONE ELSE '1';
	
	CLR_CLK_COUNT <= '0' WHEN (STATE = CS_HIGH AND CLK_COUNT = "110010") OR (STATE = CLK_HIGH AND CLK_COUNT = "110001" AND BIT_COUNT /= "10000") OR (STATE = DONE) ELSE '1';
	EN_CLK_COUNT <= '1' WHEN (STATE = CS_HIGH AND CLK_COUNT /= "110010") OR (STATE = CLK_LOW AND (CLK_COUNT /= "011000" OR CLK_COUNT = "011000")) OR
							 (STATE = CLK_HIGH AND CLK_COUNT /= "110001") ELSE '0';

	HTR_ADC_CLK <= '1' WHEN STATE = CLK_HIGH ELSE '0';
	HTR_ADC_CS <= '1' WHEN STATE = INIT OR STATE = CS_HIGH OR STATE = DONE ELSE '0';

END ARCHITECTURE BEHAVIOR;