----------------------- N bit gENeric COUNTer----------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY COUNTER IS
		GENERIC(N : INTEGER := 5);
		PORT(CLOCK		: IN STD_LOGIC;
			 RESET		: IN STD_LOGIC;
			 CLEAR  		: IN STD_LOGIC;
			 ENABLE		: IN STD_LOGIC;
			 COUNT		: BUFFER STD_LOGIC_VECTOR(N-1 DOWNTO 0)
			);
END ENTITY COUNTER;

ARCHITECTURE COUNTER of COUNTER IS 
BEGIN
	PROCESS(CLOCK,RESET)
	BEGIN
		IF(RESET = '0') THEN
			COUNT <= (OTHERS => '0');		
		ELSIF(CLOCK = '1' AND CLOCK'EVENT) THEN
			IF(CLEAR = '0') THEN
				COUNT <= (OTHERS => '0');		
			ELSIF(ENABLE = '1') THEN
				COUNT <= COUNT + 1;
			END IF;
		END IF;	
	END PROCESS;
END ARCHITECTURE COUNTER;				
---------------------------end of counter---------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY HEARTBEAT_ISA IS

PORT(CLOCK	: IN STD_LOGIC;
	  RESET	: IN STD_LOGIC;
	  	  
	  HB_ISA	: OUT STD_LOGIC
	  );
	  
END ENTITY HEARTBEAT_ISA;

ARCHITECTURE BEHAVIOR OF HEARTBEAT_ISA IS

component COUNTER IS
		GENERIC(N : INTEGER := 5);
		PORT(CLOCK		: IN STD_LOGIC;
			 RESET		: IN STD_LOGIC;
			 CLEAR  		: IN STD_LOGIC;
			 ENABLE		: IN STD_LOGIC;
			 COUNT		: BUFFER STD_LOGIC_VECTOR(N-1 DOWNTO 0)
			);
END component;

TYPE STATE_TYPE IS (S0, S1, S2, S3);
SIGNAL Y						: STATE_TYPE;

SIGNAL EN_HB_COUNT		: STD_LOGIC;
SIGNAL CLR_HB_COUNT		: STD_LOGIC;
SIGNAL HB_COUNT			: STD_LOGIC_VECTOR(26 DOWNTO 0);

BEGIN

HB_COUNTER: COUNTER
		GENERIC MAP(N => 27)
		PORT MAP(CLOCK		=> CLOCK,
					RESET		=> RESET,
					CLEAR		=> CLR_HB_COUNT,
					ENABLE	=> EN_HB_COUNT,
					COUNT		=> HB_COUNT
					);
					
	PROCESS(CLOCK, RESET)
	BEGIN
		IF RESET = '0' THEN Y <= S0;
		ELSIF (CLOCK = '1' AND CLOCK'EVENT) THEN
			CASE Y IS
			
				WHEN S0	=>	IF HB_COUNT	= "000" & X"ACFC00" THEN Y <= S1;
								ELSE Y <= S0;
								END IF;
								
				WHEN S1	=> IF HB_COUNT = "000" & X"ACFC00" THEN Y <= S2;
								ELSE Y <= S1;
								END IF;
								
				WHEN S2	=>	IF HB_COUNT = "000" & X"ACFC00" THEN Y <= S3;
								ELSE Y <= S2;
								END IF;
								
				WHEN S3	=> IF HB_COUNT = "000" & X"ACFC00" THEN Y <= S0;
								ELSE Y <= S3;
								END IF;
									
				WHEN OTHERS	=> Y <= S0;
				
			END CASE;
			
		END IF;
	END PROCESS;
		
CLR_HB_COUNT 	<= '0' WHEN ((Y = S0 OR Y = S1 OR Y = S2 OR Y = S3) AND HB_COUNT = "000" & X"ACFC00")	ELSE '1';	

EN_HB_COUNT 	<= '1' WHEN ((Y = S0 OR Y = S1 OR Y = S2 OR Y = S3) AND HB_COUNT /= "000" & X"ACFC00")	ELSE '0';


HB_ISA			<= '1' WHEN Y = S0 OR Y = S2 ELSE '0';
									

END ARCHITECTURE BEHAVIOR;