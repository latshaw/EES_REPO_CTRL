module PLL_main (
		input  wire  rst,      //   reset.reset
		input  wire  refclk,   //  refclk.clk
		output wire  outclk_0, // outclk0.clk
		output wire  outclk_1  // outclk1.clk
	);
endmodule

