LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE WORK.COMPONENTS.ALL;

ENTITY FCC_DATA_OUT IS

PORT(RESET : IN STD_LOGIC;
	  CLOCK : IN STD_LOGIC;
	  
	  RF_ON_OFF : IN STD_LOGIC;----'0'-OFF, '1'-ON
	  STEPPER_MANUAL_AUTO : IN STD_LOGIC;----'0'-MANUAL, '1'-AUTO
	  CAV_MODE : IN STD_LOGIC_VECTOR(1 DOWNTO 0);----"00"-TONE, "01"-SEL, "10"-GDR
	  
	  DISC_SMALL : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
	  DISC_MEDIUM : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
	  DISC_LARGE : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
	  DISC_XLARGE : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
	  
	  DETA : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
	  STEPS : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
	  
	  MOVE : IN STD_LOGIC;
	  DIRECTION : IN STD_LOGIC;
	  STOP : IN STD_LOGIC;
	  
	  FIBER_DATA_OUT : OUT STD_LOGIC
	  );
	  
END ENTITY FCC_DATA_OUT;

ARCHITECTURE BEHAVIOR OF FCC_DATA_OUT IS

SIGNAL FIBER_DATA_OUT_BUFFER 	: STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL EN_FIBER_DATA_OUT		: STD_LOGIC;
SIGNAL LD_FIBER_DATA_OUT		: STD_LOGIC;

SIGNAL EN_CLK_COUNT				: STD_LOGIC;
SIGNAL CLK_COUNT					: STD_LOGIC_VECTOR(2 DOWNTO 0);

SIGNAL EN_BIT_COUNT				: STD_LOGIC;
SIGNAL CLR_BIT_COUNT				: STD_LOGIC;
SIGNAL BIT_COUNT					: STD_LOGIC_VECTOR(4 DOWNTO 0);

SIGNAL EN_REG_COUNT				: STD_LOGIC;
SIGNAL REG_COUNT					: STD_LOGIC_VECTOR(2 DOWNTO 0);

SIGNAL FCC_MODE					: STD_LOGIC_VECTOR(23 DOWNTO 0);
SIGNAL COMMAND						: STD_LOGIC_VECTOR(23 DOWNTO 0);

TYPE STATE_TYPE IS (INIT, LOAD, START_TX, TX_DATA);
SIGNAL STATE						: STATE_TYPE;

BEGIN

FIBER_DATA_OUT_BUFFER(31 DOWNTO 28) <= "1000"; ------START BIT FOLLOWED BY THREE '0' BITS

-----------REGISTER STRUCTURE--------
----000-----FCC MODE(SEL, GDR, TONE, RF ON/OFF, MANUAL/AUTO)
----001-----STEPS IN THE MANUAL MODE
----010-----STEPPER COMMAND MOVE,DIRECTION,STOP
----011-----DISC SMALL
----100-----DISC MEDIUM
----101-----DISC LARGE
----110-----DISC XLARGE
----111-----DETA
FIBER_DATA_OUT_BUFFER(27 DOWNTO 25) <= REG_COUNT; -------DEFINES THE REGISTER---

FIBER_DATA_OUT_BUFFER(24 DOWNTO 1) <= STEPS WHEN REG_COUNT = "001" ELSE
												  COMMAND WHEN REG_COUNT = "010" ELSE
												  DISC_SMALL WHEN REG_COUNT = "011" ELSE
												  DISC_MEDIUM WHEN REG_COUNT = "100" ELSE
												  DISC_LARGE WHEN REG_COUNT = "101" ELSE
												  DISC_XLARGE WHEN REG_COUNT = "110" ELSE
												  DETA WHEN REG_COUNT = "111" ELSE
												  FCC_MODE;												  

FIBER_DATA_OUT_BUFFER(0) <= '0'; --------END OF TRANSMISSION BIT


COMMAND <= X"00000" & '0' & MOVE & DIRECTION & STOP;
FCC_MODE <= X"00000" & CAV_MODE & RF_ON_OFF & STEPPER_MANUAL_AUTO;

	------CLOCK COUNTER------------------------
	
	CLK_COUNTER: COUNTER
		GENERIC MAP(N => 3)
		PORT MAP(CLOCK		=> CLOCK,
					RESET		=> RESET,
					CLEAR  	=> '1',
					EN			=> EN_CLK_COUNT,
					COUNT		=> CLK_COUNT
					);
	------END OF CLOCK COUNTER------------------------
	
	------BIT COUNTER------------------------
	
	BIT_COUNTER: COUNTER
		GENERIC MAP(N => 5)
		PORT MAP(CLOCK		=> CLOCK,
					RESET		=> RESET,
					CLEAR  	=> CLR_BIT_COUNT,
					EN			=> EN_BIT_COUNT,
					COUNT		=> BIT_COUNT
					);
	------END OF BIT COUNTER------------------------


	------REGISTER COUNTER------------------------
	
	REG_COUNTER: COUNTER
		GENERIC MAP(N => 3)
		PORT MAP(CLOCK		=> CLOCK,
					RESET		=> RESET,
					CLEAR  	=> '1',
					EN			=> EN_REG_COUNT,
					COUNT		=> REG_COUNT
					);
	------END OF REGISTER COUNTER------------------------

   -------FIBER DATA OUT REGISTER----------------------
	
	FIBER_DATA_OUT_REG: SHIFT_LEFT_REG
	GENERIC MAP(N => 32)
	PORT MAP(CLOCK	=> CLOCK,
		 RESET 	=> RESET,
		 EN 		=> EN_FIBER_DATA_OUT,
		 LOAD		=> LD_FIBER_DATA_OUT,
		 CLEAR	=> '1', 
		 INP		=> FIBER_DATA_OUT_BUFFER, 
		 OUTPUT	=> FIBER_DATA_OUT 
		 );

   --------END OF FIBER DATA OUT REGISTER---------------
												  
												  
												  
												  
	PROCESS(CLOCK, RESET)
	BEGIN
		IF(RESET = '0') THEN
			STATE <= INIT;
		ELSIF(CLOCK = '1' AND CLOCK'EVENT) THEN
			
			CASE STATE IS
			
				WHEN INIT		=> STATE <= LOAD;
				
				WHEN LOAD		=> STATE <= START_TX;
				
				WHEN START_TX	=> IF(CLK_COUNT = "111") THEN STATE <= TX_DATA;
										ELSE STATE <= START_TX;
										END IF;
				
				WHEN TX_DATA	=> IF(BIT_COUNT = "11111") THEN STATE <= LOAD;
										ELSE STATE <= TX_DATA;
										END IF;
										
			END CASE;

		END IF;			
	END PROCESS;
	
EN_CLK_COUNT			<= '1' WHEN STATE = LOAD OR STATE = START_TX OR STATE = TX_DATA ELSE '0';

EN_BIT_COUNT			<= '1' WHEN (STATE = START_TX OR STATE = TX_DATA) AND (CLK_COUNT = "111") ELSE '0';
CLR_BIT_COUNT			<= '0' WHEN STATE = LOAD ELSE '1';

EN_REG_COUNT			<= '1' WHEN (STATE = TX_DATA AND BIT_COUNT = "11111") ELSE '0';

EN_FIBER_DATA_OUT 	<= '1' WHEN  (STATE = START_TX OR STATE = TX_DATA) AND (CLK_COUNT = "111") ELSE '0';
LD_FIBER_DATA_OUT		<= '1' WHEN (STATE = LOAD) ELSE '0';	


END ARCHITECTURE BEHAVIOR;
