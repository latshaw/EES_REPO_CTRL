LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE WORK.COMPONENTS.ALL;


ENTITY POLYNOMIAL_DIVISION IS
PORT(CLOCK : IN STD_LOGIC;
	  RESET : IN STD_LOGIC;
	  DATA_IN : IN STD_LOGIC_VECTOR(39 DOWNTO 0);
	  DENOM : IN STD_LOGIC_VECTOR(8 DOWNTO 0);-----x^8+x^2+x+1 ("100000111")
	  START_CRC : IN STD_LOGIC;
	  CRC : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	  DATA_OUT_CRC : OUT STD_LOGIC_VECTOR(39 DOWNTO 0);
	  CRC_DONE : OUT STD_LOGIC
	  );
END ENTITY POLYNOMIAL_DIVISION;

ARCHITECTURE BEHAVIOR OF POLYNOMIAL_DIVISION IS

SIGNAL NUMER_CRC 				: STD_LOGIC_VECTOR(39 DOWNTO 0);
SIGNAL NUMER_XOR				: STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL NUMER_CRC_REG			: STD_LOGIC_VECTOR(39 DOWNTO 0);
SIGNAL CRC_COMPARE			: STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL NUMER_CRC_BIT			: STD_LOGIC;

SIGNAL EN_CRC_REG				: STD_LOGIC;
SIGNAL LD_CRC_REG				: STD_LOGIC;

SIGNAL CRC_INPUT				: STD_LOGIC_VECTOR(7 DOWNTO 0);

SIGNAL EN_CRC_RESULT			: STD_LOGIC;

SIGNAL EN_DATA					: STD_LOGIC;

SIGNAL CLR_SHIFT_COUNT		: STD_LOGIC;
SIGNAL EN_SHIFT_COUNT		: STD_LOGIC;
SIGNAL SHIFT_COUNT			: STD_LOGIC_VECTOR(4 DOWNTO 0);

SIGNAL EN_XOR_SHIFT			: STD_LOGIC;
SIGNAL LD_XOR_SHIFT			: STD_LOGIC;
SIGNAL INP_XOR_SHIFT			: STD_LOGIC_VECTOR(8 DOWNTO 0);
SIGNAL OUP_XOR_SHIFT			: STD_LOGIC_VECTOR(8 DOWNTO 0);

SIGNAL INP_XOR_SHIFT_SEL	: STD_LOGIC_VECTOR(8 DOWNTO 0);

SIGNAL SHIFT_SEL				: STD_LOGIC;

SIGNAL EN_DATA_OUT			: STD_LOGIC;
SIGNAL DATA_OUT				: STD_LOGIC_VECTOR(39 DOWNTO 0);

SIGNAL CRC_DONE_TMP			: STD_LOGIC;


TYPE STATE_TYPE IS (INIT, LOAD_NUMER, LOAD_NUMER_WAIT, LOAD_XOR_INIT, EN_XOR, CHECK_MSB, EN_NUMER, LOAD_XOR, RESULT);
SIGNAL STATE					: STATE_TYPE;

BEGIN

NUMER_CRC <= DATA_IN;


DATA_OUT <= NUMER_CRC_REG (39 DOWNTO 8)& OUP_XOR_SHIFT(7 DOWNTO 0);

INP_XOR_SHIFT <= INP_XOR_SHIFT_SEL XOR DENOM;

INP_XOR_SHIFT_SEL <=  OUP_XOR_SHIFT WHEN SHIFT_SEL = '1' ELSE  NUMER_CRC_REG(39 DOWNTO 31);

--------------------CRC_DONE_OUT FLIP FLOP-------------------


CRC_DONE_FF: LATCH_N 
	PORT MAP(CLOCK	=> CLOCK, 
				RESET => RESET,
				CLEAR => '1', 
				EN 	=> '1',
				INP 	=> CRC_DONE_TMP,
				OUP	=> CRC_DONE 
				);

---------------REGISTER FOR THE DATA TO BE PROCESSED FOR CRC------------------------
NUMER_REG: REGNE
		GENERIC MAP(N => 40) 
		PORT MAP(CLOCK		=> CLOCK,
					RESET 	=> RESET,
					CLEAR		=> '1',  
					EN			=> EN_DATA,
					INPUT		=> NUMER_CRC,
					OUTPUT	=> NUMER_CRC_REG
					);
					
---------------REGISTER FOR DATA OUT------------------------
DATA_OUT_REG: REGNE
		GENERIC MAP(N => 40) 
		PORT MAP(CLOCK		=> CLOCK,
					RESET 	=> RESET,
					CLEAR		=> '1',  
					EN			=> EN_DATA_OUT,
					INPUT		=> DATA_OUT,
					OUTPUT	=> DATA_OUT_CRC
					);


-------REGISTER FOR 31 BITS THAT WILL BE SHIFTED FOR CALCULATING CRC-----------------
					
NUMER_CRC_SHIFT_REG: SHIFT_LEFT_REG
	GENERIC MAP(N => 31)
	PORT MAP(CLOCK		=> CLOCK,	
				RESET		=> RESET,
				EN			=> EN_CRC_REG,
				CLEAR		=> '1',
				LOAD		=> LD_CRC_REG,
				INP		=> NUMER_CRC_REG(30 DOWNTO 0),
				OUTPUT	=> NUMER_CRC_BIT
				);			
				
----------REGISTER FOR 9 BIT REGISTER (XOR AND SHIFT INPUT BIT FROM NUMERATOR)----------------
				
XOR_SHIFT_REG: SHIFT_LEFT_BIT
	GENERIC MAP(N => 9)
	PORT MAP(CLOCK			=> CLOCK,	
				RESET			=> RESET,
				EN				=> EN_XOR_SHIFT,
				LOAD			=> LD_XOR_SHIFT,
				SHIFT_BIT	=> NUMER_CRC_BIT,
				INP			=> INP_XOR_SHIFT,
				OUTPUT		=> OUP_XOR_SHIFT
				);				
				
CRC_RESULT_REG: REGNE
		GENERIC MAP(N => 8) 
		PORT MAP(CLOCK		=> CLOCK,
					RESET 	=> RESET,
					CLEAR		=> '1',  
					EN			=> EN_CRC_RESULT,
					INPUT		=> OUP_XOR_SHIFT(7 DOWNTO 0),
					OUTPUT	=> CRC
					);
					
SHIFT_BIT_COUNTER: COUNTER
		GENERIC MAP(N => 5)
		PORT MAP(CLOCK		=> CLOCK,	
					RESET		=> RESET,
					CLEAR		=> CLR_SHIFT_COUNT,
					EN			=> EN_SHIFT_COUNT,
					COUNT		=> SHIFT_COUNT
					);
					
					
					
	PROCESS(CLOCK, RESET)
	BEGIN
		IF(RESET = '0') THEN
			STATE <= INIT;
		ELSIF (CLOCK = '1' AND CLOCK'EVENT) THEN
			
			CASE STATE IS
				
				WHEN INIT				=> IF START_CRC = '1' THEN STATE <= LOAD_NUMER;
												ELSE STATE <= INIT;
												END IF;
												
				WHEN LOAD_NUMER		=> STATE <= LOAD_NUMER_WAIT;
				
				WHEN LOAD_NUMER_WAIT	=> STATE <= LOAD_XOR_INIT;
									
				WHEN LOAD_XOR_INIT	=> STATE <= EN_XOR;
				
				WHEN EN_XOR				=> STATE <= CHECK_MSB;
				
				
				WHEN CHECK_MSB			=> IF OUP_XOR_SHIFT(8) = '0' THEN
													IF SHIFT_COUNT = "11110" THEN STATE <= RESULT;
													ELSE STATE <= EN_NUMER;
													END IF;
												ELSE STATE <= LOAD_XOR;
												END IF;
												
				WHEN LOAD_XOR			=> IF SHIFT_COUNT = "11110" THEN STATE <= RESULT;
												ELSE STATE <= EN_NUMER;
												END IF;
												
				WHEN EN_NUMER			=> STATE <= EN_XOR;
		
										
				WHEN RESULT				=> STATE <= INIT;
				
				WHEN OTHERS				=> STATE <= INIT;
				
			END CASE;
		END IF;
	END PROCESS;
	
LD_CRC_REG <= '1' WHEN STATE = LOAD_NUMER_WAIT ELSE '0';
EN_CRC_REG <= '1' WHEN STATE = EN_NUMER ELSE '0';
	
EN_DATA <= '1' WHEN STATE = LOAD_NUMER ELSE '0';

EN_DATA_OUT <= '1' WHEN STATE = RESULT ELSE '0';

SHIFT_SEL <= '0' WHEN STATE = LOAD_NUMER OR STATE = LOAD_XOR_INIT ELSE '1';
		
EN_CRC_RESULT <= '1' WHEN STATE = RESULT ELSE '0';
					
EN_XOR_SHIFT <= '1' WHEN STATE = EN_XOR ELSE '0';

LD_XOR_SHIFT <= '1' WHEN STATE = LOAD_XOR_INIT OR STATE = LOAD_XOR ELSE '0';

EN_SHIFT_COUNT <= '1' WHEN STATE = EN_NUMER ELSE '0';
CLR_SHIFT_COUNT <= '0' WHEN STATE = LOAD_NUMER ELSE '1';

CRC_DONE_TMP <= '1' WHEN STATE = RESULT ELSE '0';

END ARCHITECTURE BEHAVIOR;