--LIBRARY IEEE;
--USE IEEE.STD_LOGIC_1164.ALL;
--USE IEEE.STD_LOGIC_UNSIGNED.ALL;
--USE WORK.COMPONENTS.ALL;
--
--ENTITY IIR_SIMPLE IS
--
--PORT(RESET 	: IN STD_LOGIC;
--	 CLOCK 	: IN STD_LOGIC;
--	 LOAD	: IN STD_LOGIC;
--	 I		: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
--	 O		: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
--	 );
--	  
--END ENTITY IIR_SIMPLE;
--
--ARCHITECTURE BEHAVIOR OF IIR_SIMPLE IS
--
--SIGNAL I_EXT		: STD_LOGIC_VECTOR(36 DOWNTO 0);
--SIGNAL REG_SHIFT	: STD_LOGIC_VECTOR(36 DOWNTO 0);
--SIGNAL REG			: STD_LOGIC_VECTOR(36 DOWNTO 0);
--
--SIGNAL ONE			: STD_LOGIC;
--
--SIGNAL REG_IN		: STD_LOGIC_VECTOR(36 DOWNTO 0);
--SIGNAL REG_OUT		: STD_LOGIC_VECTOR(36 DOWNTO 0);
--
--
--
--BEGIN
--
--ONE <= '1';
--
--
--
---- extend the input to 32 bits
--I_EXT(36 DOWNTO 16) <= (OTHERS => I(15));
--I_EXT(15 DOWNTO 0)  <= I;
--
---- setup register
--FILTER_REG: REGNE
--		GENERIC MAP(N => 37) 
--		PORT MAP(CLOCK		=> CLOCK,
--					RESET		=> RESET,
--					CLEAR		=> ONE,
--					EN			=> LOAD,	
--					INPUT		=> REG_IN,
--					OUTPUT	=> REG_OUT
--					);
--					
--
--
--					
--REG_IN <= REG_OUT + I_EXT - REG_SHIFT;
--
--
--
--			REG_SHIFT(36 DOWNTO 17) <= (OTHERS => REG_OUT(36));
--			REG_SHIFT(16 DOWNTO 0)  <= REG_OUT(36 DOWNTO 20);
--			
--			
--			O <= REG_IN(35 DOWNTO 20) WHEN REG_IN(36 DOWNTO 35) = "00" OR REG_IN(36 DOWNTO 35) = "11" ELSE
--				  X"7FFF" WHEN REG_IN(36 DOWNTO 35) = "01" ELSE
--				  X"8000";
--				  
--END ARCHITECTURE BEHAVIOR;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE WORK.COMPONENTS.ALL;

ENTITY IIR_SIMPLE IS

PORT(CLOCK 	: IN STD_LOGIC;
	  RESET 	: IN STD_LOGIC;
	  LOAD	: IN STD_LOGIC;
	  I		: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	  O		: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	  );
	  
END ENTITY IIR_SIMPLE;

ARCHITECTURE BEHAVIOR OF IIR_SIMPLE IS

SIGNAL I_EXT		: STD_LOGIC_VECTOR(33 DOWNTO 0);
SIGNAL REG_SHIFT	: STD_LOGIC_VECTOR(33 DOWNTO 0);
SIGNAL REG			: STD_LOGIC_VECTOR(33 DOWNTO 0);

SIGNAL ONE			: STD_LOGIC;

SIGNAL REG_IN		: STD_LOGIC_VECTOR(33 DOWNTO 0);
SIGNAL REG_OUT		: STD_LOGIC_VECTOR(33 DOWNTO 0);

SIGNAL O_INT		: STD_LOGIC_VECTOR(15 DOWNTO 0);



BEGIN

ONE <= '1';



-- extend the input to 30 bits
I_EXT(33 DOWNTO 16) <= (OTHERS => I(15));
I_EXT(15 DOWNTO 0)  <= I;

-- setup register
FILTER_REG: REGNE
		GENERIC MAP(N => 34) 
		PORT MAP(CLOCK		=> CLOCK,
					RESET		=> RESET,
					CLEAR		=> ONE,
					EN			=> LOAD,	
					INPUT		=> REG_IN,
					OUTPUT	=> REG_OUT
					);
					


					
REG_IN <= REG_OUT - REG_SHIFT + I_EXT;



			REG_SHIFT(33 DOWNTO 24) <= (OTHERS => REG_OUT(33));
			REG_SHIFT(23 DOWNTO 0)  <= REG_OUT(33 DOWNTO 10);
			
			
			O_INT <= X"7FFF" WHEN REG_OUT(33) = '0' AND REG_OUT(32 DOWNTO 25) /= ("00000000") ELSE
				  X"8000" WHEN REG_OUT(33) = '1' AND REG_OUT(32 DOWNTO 25) /= ("11111111") ELSE
				  REG_OUT(25 DOWNTO 10);
				  
OUTPUT_REG: REGNE
		GENERIC MAP(N => 16) 
		PORT MAP(CLOCK		=> CLOCK,
					RESET		=> RESET,
					CLEAR		=> ONE,
					EN			=> LOAD,	
					INPUT		=> O_INT,
					OUTPUT	=> O
					);
				  
END ARCHITECTURE BEHAVIOR;