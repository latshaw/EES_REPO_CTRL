LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE WORK.COMPONENTS.ALL;

ENTITY DATA_SELECT IS

PORT(STEPS_FIB : IN REG32_ARRAY;     
	  DIR_FIB : IN STD_LOGIC_VECTOR(7 DOWNTO 0);	  
	  MOVE_FIB : IN STD_LOGIC_VECTOR(7 DOWNTO 0);	  
	  DONE_FIB : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  FIB_MODE : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  
	  STEPS : IN REG32_ARRAY;	  
	  DIR : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  MOVE : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  DONE : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	  
	  STEPS_OUT : OUT REG32_ARRAY;
	  DIR_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	  MOVE_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	  DONE_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	  );
	  
END ENTITY DATA_SELECT;

ARCHITECTURE BEHAVIOR OF DATA_SELECT IS

SIGNAL DONE_FIB_CHK	: STD_LOGIC_VECTOR(7 DOWNTO 0);

BEGIN

DATA_MUX_GEN: FOR I IN 0 TO 7 GENERATE


DONE_FIB_CHK(I) <= '0' WHEN (STEPS_FIB(I) = x"00000000") ELSE DONE_FIB(I);

DONE_OUT(I) <= DONE_FIB_CHK(I) WHEN FIB_MODE(I) = '1' ELSE DONE(I);
STEPS_OUT(I)(31 DOWNTO 0) <= STEPS_FIB(I)(31 DOWNTO 0) WHEN FIB_MODE(I) = '1' ELSE STEPS(I)(31 DOWNTO 0);
DIR_OUT(I) <= DIR_FIB(I) WHEN FIB_MODE(I) = '1' ELSE DIR(I);
MOVE_OUT(I) <= MOVE_FIB(I) WHEN FIB_MODE(I) = '1' ELSE MOVE(I);

END GENERATE;

END ARCHITECTURE BEHAVIOR;
	  