-- llrf 3.0 note, i am adding comments to this module to understand how it worked, however we will be using
-- the ads8353 adc in place of this adc so the f/w will be different.

-- this moduel contols 2, 4 channel adc (8 analog values being digitized)

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE WORK.COMPONENTS.ALL;

ENTITY AD7367_CONTROL IS

PORT(CLOCK : IN STD_LOGIC;
	 RESET : IN STD_LOGIC;
	 ARC_ADC_BSY : IN STD_LOGIC;
	 ARC_ADC1_DOUTA : IN STD_LOGIC;
	 ARC_ADC1_DOUTB : IN STD_LOGIC;
	 ARC_ADC2_DOUTA : IN STD_LOGIC;
	 ARC_ADC2_DOUTB : IN STD_LOGIC;
	 ARC_TRIG_DELAY : IN REG16_ARRAY;
	 ARC_STOP : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	 ARC_FAULT_CLEAR : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	 ARC_FAULT : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	 ARC_BUF_ADDR_IN : IN STD_LOGIC_VECTOR(15 DOWNTO 1);
	 
	 ARC_DATA : OUT REG16_ARRAY; -- outputs arc data value, channel specific
	 
	 ARC_BUF_EN : OUT STD_LOGIC_VECTOR(7 DOWNTO 0); -- these buffer address are not clear to me. ARC_BUF_ADDR is either the adc write address or the adc read address (after stop or fault is hi for the specified number of deay ticks)
	 ARC_BUF_ADDR : OUT REG11_ARRAY;
	 ARC_ADC_CNVST : OUT STD_LOGIC;
	 ARC_ADC_CS : OUT STD_LOGIC;
	 ARC_ADC_SCLK : OUT STD_LOGIC;
	 ARC_ADC_ADDR : OUT STD_LOGIC;
	 ARC_BUFF_READY : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	 
	 --COMPARE : OUT STD_LOGIC;
	 
	 --DAC_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	 
	 );
END ENTITY AD7367_CONTROL;

ARCHITECTURE BEHAVIOR OF AD7367_CONTROL IS


SIGNAL ARC_ADC_ADDR_TEMP	: STD_LOGIC_VECTOR(1 DOWNTO 0);

SIGNAL SCLK_COUNT			: STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL EN_SCLK_COUNT		: STD_LOGIC;
SIGNAL CLEAR_SCLK_COUNT		: STD_LOGIC;

SIGNAL BIT_COUNT			: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL EN_BIT_COUNT			: STD_LOGIC;
SIGNAL CLEAR_BIT_COUNT		: STD_LOGIC;

SIGNAL EN_DOUT				: STD_LOGIC;

SIGNAL CLEAR_ARC_COUNT		: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL EN_ARC_BUF_COUNT		: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL ARC_WRITE_ADDR		: REG11_ARRAY;

SIGNAL ARC_DATA_IN			: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL ARC_DATA_TEMP		: REG14_ARRAY;
SIGNAL ARC_DATA_REG_IN		: REG16_ARRAY;
SIGNAL EN_ARC_DATA_REG		: STD_LOGIC;
SIGNAL EN_ARC_DATA			: STD_LOGIC_VECTOR(7 DOWNTO 0);

SIGNAL EN_ARC_ADDR			: STD_LOGIC;

SIGNAL CLR_ARC_ADDR			: STD_LOGIC;

SIGNAL ARC_READ_ADDR		: REG12_ARRAY;

SIGNAL ARC_READ_LATCH_ADDR	: REG11_ARRAY;


signal ONE					: STD_LOGIC;

SIGNAL CLR_ARC_TRIG_COUNT	: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL EN_ARC_TRIG_COUNT	: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL ARC_TRIG_COUNT		: REG16_ARRAY;
SIGNAL ARC_TRIG_DONE		: STD_LOGIC_VECTOR(7 DOWNTO 0);

SIGNAL ARC_FAULT_STOP		: STD_LOGIC_VECTOR(7 DOWNTO 0);

SIGNAL ARC_BUF_DIS			: STD_LOGIC_VECTOR(7 DOWNTO 0);

TYPE STATE_TYPE IS (INIT, CONVERT, BUSY, ACQUIRE, CS_WAIT, SCLK_LOW, SCLK_HIGH, T_QUIET);
SIGNAL STATE : STATE_TYPE;

attribute ENUM_ENCODING: STRING;

attribute ENUM_ENCODING of STATE_TYPE:type is "00000001 00000010 00000100 00001000 00010000 00100000 01000000 10000000" ;

BEGIN

ONE <= '1';
--arc_trig_test <= x"03e8";

-----ARC TRIGGER DELAY COUNTERS-----------------

ARC_TRIG_CNT_GEN: FOR I IN 0 TO 7 GENERATE
	-- counter to ensure that the channel specific number of ARC_TRIG_DELAY ticks/counts have occured
	ARC_TRIG_COUNTERI: COUNTER
		GENERIC MAP(N => 16)
		PORT MAP(CLOCK	=> CLOCK,	
				 RESET	=> RESET,
				 CLEAR  => NOT ARC_FAULT_CLEAR(I),--CLR_ARC_TRIG_COUNT(I),
				 ENABLE	=> EN_ARC_TRIG_COUNT(I),
				 COUNT	=> ARC_TRIG_COUNT(I)
				);
			

	-- enable counter when either arc fault or arc stop input are hi
	EN_ARC_TRIG_COUNT(I) <= '1' WHEN (ARC_FAULT_STOP(I) = '1' AND ARC_TRIG_DONE(I) = '0') ELSE '0';
	
	-- trigger counter has completed
	ARC_TRIG_DONE(I) <= '1' WHEN ARC_TRIG_COUNT(I) = ARC_TRIG_DELAY(I) ELSE '0';---commented out for testing
	
	--arc buffer display
	ARC_BUF_DIS(I) <= '1' WHEN (ARC_FAULT_STOP(I) = '1' AND ARC_TRIG_DONE(I) = '1') ELSE '0'; --buffer write is disabled when arc stop or arc fault occurs
																															--and samples are taken for trig delay after the fault					
	-- will go hi if the module has an arc fault input or an arc stop input
	ARC_FAULT_STOP(I) <= ARC_FAULT(I) OR ARC_STOP(I);										  
			
END GENERATE;

-- channel specific signal, when this is HI, it means that the ARC_FAULT(I) OR ARC_STOP(I) have been hi for ARC_TRIG_DELAY number of ticks
ARC_BUFF_READY <= ARC_TRIG_DONE;

--------------------------------------------------

GEN_REG_ARC: FOR I IN 0 TO 7 GENERATE	
	-- when address is selected, begin to shift in data
	SHIFT_REG_ARCI: SHIFT_LEFT_REG
		GENERIC MAP(N => 14)
		PORT MAP(CLOCK	=> CLOCK, 
				 RESET	=> RESET,
				 EN		=> EN_ARC_DATA(I),
				 INP	=> ARC_DATA_IN(I),
				 OUTPUT	=> ARC_DATA_TEMP(I)
				);
					
				
	ARC_DATA_REG: REGNE
		GENERIC MAP(N => 16) 
		PORT MAP(CLOCK 	=> CLOCK,
				 RESET 	=> RESET,
				 CLEAR  => ONE,
				 EN		=> EN_ARC_DATA_REG,
				 INPUT	=> ARC_DATA_REG_IN(I),
				 OUTPUT => ARC_DATA(I) -- holds the registered arc data value, module output
				);
	-- place holder for data being shifted in 			
	ARC_DATA_REG_IN(I) 		<= "00" & NOT ARC_DATA_TEMP(I)(13) & ARC_DATA_TEMP(I)(12 DOWNTO 0);
	
END GENERATE;
	-- when this is hi, data is ready to be registered (done shifitng in data for that line)
	EN_ARC_DATA_REG 		<= '1' WHEN (STATE = SCLK_LOW AND BIT_COUNT = "1101" AND SCLK_COUNT = "10") ELSE '0';
	
	
ARC_ADDR_GEN: FOR I IN 0 TO 7 GENERATE
	
	ARC_WRITE_ADDR_COUNTERI: COUNTER
		GENERIC MAP(N => 11)
		PORT MAP(CLOCK	=> CLOCK,	
			 RESET	=> RESET,
			 CLEAR  => ONE,--CLEAR_ARC_COUNT(I),
			 ENABLE	=> EN_ARC_BUF_COUNT(I),
			 COUNT	=> ARC_WRITE_ADDR(I)
			);
			
	

	--ARC_BUF_ADDR(I) <= arc_write_addr(i);---for testing
			
	--CLEAR_ARC_COUNT(I) <= ONE;
			
END GENERATE;


-- 						
ARC_BUF_ADDR(0) <= ARC_READ_ADDR(0)(10 DOWNTO 0) WHEN (ARC_BUF_DIS(0) = '1' AND ARC_BUF_ADDR_IN(15 DOWNTO 12) = x"4") ELSE ARC_WRITE_ADDR(0);---commented out for testing
ARC_BUF_ADDR(1) <= ARC_READ_ADDR(1)(10 DOWNTO 0) WHEN (ARC_BUF_DIS(1) = '1' AND ARC_BUF_ADDR_IN(15 DOWNTO 12) = x"5") ELSE ARC_WRITE_ADDR(1);
ARC_BUF_ADDR(2) <= ARC_READ_ADDR(2)(10 DOWNTO 0) WHEN (ARC_BUF_DIS(2) = '1' AND ARC_BUF_ADDR_IN(15 DOWNTO 12) = x"6") ELSE ARC_WRITE_ADDR(2);
ARC_BUF_ADDR(3) <= ARC_READ_ADDR(3)(10 DOWNTO 0) WHEN (ARC_BUF_DIS(3) = '1' AND ARC_BUF_ADDR_IN(15 DOWNTO 12) = x"7") ELSE ARC_WRITE_ADDR(3);
ARC_BUF_ADDR(4) <= ARC_READ_ADDR(4)(10 DOWNTO 0) WHEN (ARC_BUF_DIS(4) = '1' AND ARC_BUF_ADDR_IN(15 DOWNTO 12) = x"8") ELSE ARC_WRITE_ADDR(4);
ARC_BUF_ADDR(5) <= ARC_READ_ADDR(5)(10 DOWNTO 0) WHEN (ARC_BUF_DIS(5) = '1' AND ARC_BUF_ADDR_IN(15 DOWNTO 12) = x"9") ELSE ARC_WRITE_ADDR(5);
ARC_BUF_ADDR(6) <= ARC_READ_ADDR(6)(10 DOWNTO 0) WHEN (ARC_BUF_DIS(6) = '1' AND ARC_BUF_ADDR_IN(15 DOWNTO 12) = x"A") ELSE ARC_WRITE_ADDR(6);
ARC_BUF_ADDR(7) <= ARC_READ_ADDR(7)(10 DOWNTO 0) WHEN (ARC_BUF_DIS(7) = '1' AND ARC_BUF_ADDR_IN(15 DOWNTO 12) = x"B") ELSE ARC_WRITE_ADDR(7);








ARC_BUF_READ_ADDR_GEN: FOR I IN 0 TO 7 GENERATE----- REGISTERTING THE ADDRESS WHEN BUFFER IS DISABLED
											----- WHEN ARC_STOP_BUF IS '1' AND ARC_TRIG_DONE = '1'
	ARC_BUF_READ_ADDR_GEN: REGNE
		GENERIC MAP(N => 11) 
		PORT MAP(CLOCK 	=> CLOCK,
				 RESET 	=> RESET,
				 CLEAR  => ONE,
				 EN		=> ARC_TRIG_DONE(I),
				 INPUT	=> ARC_WRITE_ADDR(I),
				 OUTPUT => ARC_READ_LATCH_ADDR(I)----THIS IS THE MOST RECENT SAMPLE
				);
				
-----DEFINING ARC_READ_ADDR BASED ON ARC_READ_LATCH_ADDR AND INCOMING ISA READ ADDRESS
	ARC_READ_ADDR(I) <= ('0' & ARC_READ_LATCH_ADDR(I)) + ARC_BUF_ADDR_IN(11 DOWNTO 1) + '1';----ADDING '1' TO POINT TO THE OLDEST SAMPLE
				
END GENERATE;

	EN_ARC_BUF_COUNT(0) <= '1' WHEN (STATE = T_QUIET AND BIT_COUNT = "1110" AND ARC_ADC_ADDR_TEMP(0) = '1' AND ARC_BUF_DIS(0) = '0') ELSE '0';
	EN_ARC_BUF_COUNT(1) <= '1' WHEN (STATE = T_QUIET AND BIT_COUNT = "1110" AND ARC_ADC_ADDR_TEMP(0) = '0' AND ARC_BUF_DIS(1) = '0') ELSE '0';
	EN_ARC_BUF_COUNT(2) <= '1' WHEN (STATE = T_QUIET AND BIT_COUNT = "1110" AND ARC_ADC_ADDR_TEMP(0) = '0' AND ARC_BUF_DIS(2) = '0') ELSE '0';
	EN_ARC_BUF_COUNT(3) <= '1' WHEN (STATE = T_QUIET AND BIT_COUNT = "1110" AND ARC_ADC_ADDR_TEMP(0) = '1' AND ARC_BUF_DIS(3) = '0') ELSE '0';
	EN_ARC_BUF_COUNT(4) <= '1' WHEN (STATE = T_QUIET AND BIT_COUNT = "1110" AND ARC_ADC_ADDR_TEMP(0) = '1' AND ARC_BUF_DIS(4) = '0') ELSE '0';
	EN_ARC_BUF_COUNT(5) <= '1' WHEN (STATE = T_QUIET AND BIT_COUNT = "1110" AND ARC_ADC_ADDR_TEMP(0) = '0' AND ARC_BUF_DIS(5) = '0') ELSE '0';
	EN_ARC_BUF_COUNT(6) <= '1' WHEN (STATE = T_QUIET AND BIT_COUNT = "1110" AND ARC_ADC_ADDR_TEMP(0) = '0' AND ARC_BUF_DIS(6) = '0') ELSE '0';
	EN_ARC_BUF_COUNT(7) <= '1' WHEN (STATE = T_QUIET AND BIT_COUNT = "1110" AND ARC_ADC_ADDR_TEMP(0) = '1' AND ARC_BUF_DIS(7) = '0') ELSE '0';

	ARC_BUF_EN(0) <= '1' WHEN (STATE = SCLK_LOW AND BIT_COUNT = "1101" AND SCLK_COUNT = "11" AND ARC_ADC_ADDR_TEMP(0) = '1' AND ARC_BUF_DIS(0) = '0') ELSE '0';
	ARC_BUF_EN(1) <= '1' WHEN (STATE = SCLK_LOW AND BIT_COUNT = "1101" AND SCLK_COUNT = "11" AND ARC_ADC_ADDR_TEMP(0) = '0' AND ARC_BUF_DIS(1) = '0') ELSE '0';
	ARC_BUF_EN(2) <= '1' WHEN (STATE = SCLK_LOW AND BIT_COUNT = "1101" AND SCLK_COUNT = "11" AND ARC_ADC_ADDR_TEMP(0) = '0' AND ARC_BUF_DIS(2) = '0') ELSE '0';
	ARC_BUF_EN(3) <= '1' WHEN (STATE = SCLK_LOW AND BIT_COUNT = "1101" AND SCLK_COUNT = "11" AND ARC_ADC_ADDR_TEMP(0) = '1' AND ARC_BUF_DIS(3) = '0') ELSE '0';
	ARC_BUF_EN(4) <= '1' WHEN (STATE = SCLK_LOW AND BIT_COUNT = "1101" AND SCLK_COUNT = "11" AND ARC_ADC_ADDR_TEMP(0) = '1' AND ARC_BUF_DIS(4) = '0') ELSE '0';
	ARC_BUF_EN(5) <= '1' WHEN (STATE = SCLK_LOW AND BIT_COUNT = "1101" AND SCLK_COUNT = "11" AND ARC_ADC_ADDR_TEMP(0) = '0' AND ARC_BUF_DIS(5) = '0') ELSE '0';
	ARC_BUF_EN(6) <= '1' WHEN (STATE = SCLK_LOW AND BIT_COUNT = "1101" AND SCLK_COUNT = "11" AND ARC_ADC_ADDR_TEMP(0) = '0' AND ARC_BUF_DIS(6) = '0') ELSE '0';
	ARC_BUF_EN(7) <= '1' WHEN (STATE = SCLK_LOW AND BIT_COUNT = "1101" AND SCLK_COUNT = "11" AND ARC_ADC_ADDR_TEMP(0) = '1' AND ARC_BUF_DIS(7) = '0') ELSE '0';



	-- mapping each analog input to its respective SDO line (note, there are two, four channel adcs = 8 channels in total)
	ARC_DATA_IN(0) <= ARC_ADC1_DOUTB;--CORRESPONDS TO CAVITY 1
	ARC_DATA_IN(1) <= ARC_ADC1_DOUTB;--CORRESPONDS TO CAVITY 2
	ARC_DATA_IN(2) <= ARC_ADC1_DOUTA;--CORRESPONDS TO CAVITY 3
	ARC_DATA_IN(3) <= ARC_ADC1_DOUTA;--CORRESPONDS TO CAVITY 4 
	ARC_DATA_IN(4) <= ARC_ADC2_DOUTB;--CORRESPONDS TO CAVITY 5
	ARC_DATA_IN(5) <= ARC_ADC2_DOUTB;--CORRESPONDS TO CAVITY 6
	ARC_DATA_IN(6) <= ARC_ADC2_DOUTA;--CORRESPONDS TO CAVITY 7
	ARC_DATA_IN(7) <= ARC_ADC2_DOUTA;--CORRESPONDS TO CAVITY 8

	-- use the above adc_data_in line whenever the state machine has the correct address selected
	-- for each SDO_A and SDO_B, there are two analog channels
	EN_ARC_DATA(0) <= '1' WHEN EN_DOUT = '1' AND (ARC_ADC_ADDR_TEMP(0) = '1') ELSE '0';--CORRESPONDS TO CAVITY 1
	EN_ARC_DATA(1) <= '1' WHEN EN_DOUT = '1' AND (ARC_ADC_ADDR_TEMP(0) = '0') ELSE '0';--CORRESPONDS TO CAVITY 2
	EN_ARC_DATA(2) <= '1' WHEN EN_DOUT = '1' AND (ARC_ADC_ADDR_TEMP(0) = '0') ELSE '0';--CORRESPONDS TO CAVITY 3
	EN_ARC_DATA(3) <= '1' WHEN EN_DOUT = '1' AND (ARC_ADC_ADDR_TEMP(0) = '1') ELSE '0';--CORRESPONDS TO CAVITY 4
	EN_ARC_DATA(4) <= '1' WHEN EN_DOUT = '1' AND (ARC_ADC_ADDR_TEMP(0) = '1') ELSE '0';--CORRESPONDS TO CAVITY 5
	EN_ARC_DATA(5) <= '1' WHEN EN_DOUT = '1' AND (ARC_ADC_ADDR_TEMP(0) = '0') ELSE '0';--CORRESPONDS TO CAVITY 6
	EN_ARC_DATA(6) <= '1' WHEN EN_DOUT = '1' AND (ARC_ADC_ADDR_TEMP(0) = '0') ELSE '0';--CORRESPONDS TO CAVITY 7
	EN_ARC_DATA(7) <= '1' WHEN EN_DOUT = '1' AND (ARC_ADC_ADDR_TEMP(0) = '1') ELSE '0';--CORRESPONDS TO CAVITY 8


-- below looks like spi state machine, configures, steps through address, and extractes sdo bits


	SCLK_COUNTER: COUNTER
		GENERIC MAP(N => 2)
		PORT MAP(CLOCK	=> CLOCK,	
			 RESET	=> RESET,
			 CLEAR  => CLEAR_SCLK_COUNT,
			 ENABLE	=> EN_SCLK_COUNT,
			 COUNT	=> SCLK_COUNT
			);
			
	BIT_COUNTER: COUNTER
		GENERIC MAP(N => 4)
		PORT MAP(CLOCK	=> CLOCK,	
			 RESET	=> RESET,
			 CLEAR  => CLEAR_BIT_COUNT,
			 ENABLE	=> EN_BIT_COUNT,
			 COUNT	=> BIT_COUNT
			);
			

	ARC_ADC_COUNT: COUNTER
		GENERIC MAP(N => 2)
		PORT MAP(CLOCK => CLOCK, 
				 RESET => RESET,
				 CLEAR => CLR_ARC_ADDR,
				 ENABLE => EN_ARC_ADDR,
				 COUNT => ARC_ADC_ADDR_TEMP
				);			
			
			
	ARC_ADC_ADDR <= ARC_ADC_ADDR_TEMP(0);



	PROCESS(CLOCK, RESET, ARC_ADC_BSY, SCLK_COUNT, BIT_COUNT)
	BEGIN
		IF(RESET = '0') THEN
			STATE <= INIT;
		ELSIF(CLOCK = '1' AND CLOCK'EVENT) THEN
		
			CASE STATE IS
				
				WHEN INIT		=>	STATE <= CONVERT;		
				
				WHEN CONVERT	=>	 -- MAKING CNVST SIGNAL LOW FOR ONE CLOCK CYCLE
									IF(ARC_ADC_BSY = '0') THEN STATE <= CONVERT;
									ELSE STATE <= BUSY;
									END IF;
									
				WHEN BUSY		=>	
									IF(ARC_ADC_BSY = '1') THEN STATE <= BUSY; -- WAITING FOR BUSY SIGNAL TO GO LOW
									ELSE STATE <= ACQUIRE;
									END IF;
									
				WHEN ACQUIRE	=>	 -- MAKING CS SIGNAL LOW FOR READING THE DATA
									STATE <= CS_WAIT;
									
				
									
				WHEN CS_WAIT	=>	 
										STATE <= SCLK_HIGH;
										
										
				
				WHEN SCLK_HIGH	=>	
									
									 -- MAKING SCLK HIGH FOR 2 CLOCK CYCLES(50nS, 20 MHz)
									IF(SCLK_COUNT = "01") THEN										
										STATE <= SCLK_LOW;
									ELSE										
										STATE <= SCLK_HIGH;
									END IF;
									
				WHEN SCLK_LOW	=>	 -- MAKING SCLK LOW FOR 2 CLOCK CYCLES
									IF(SCLK_COUNT = "11") THEN
										IF(BIT_COUNT = "1101") THEN STATE <= T_QUIET;
										ELSE STATE <= SCLK_HIGH;
										END IF;
									ELSE								
										STATE <= SCLK_LOW;
									END IF;
										 
				WHEN T_QUIET	=>	
									IF(BIT_COUNT = "1111") THEN -- WAITING FOR 4 CLOCK CYCLES (T-QUIET) BEFORE NEXT CONVERSION										
										STATE <= CONVERT;
									ELSE										
										STATE <= T_QUIET;
									END IF;
								
				WHEN OTHERS		=> STATE <= INIT;	
									
			END CASE;
		END IF;
	END PROCESS;
	
	
	ARC_ADC_CNVST <= '0' WHEN STATE = CONVERT ELSE '1';
	ARC_ADC_SCLK <= '0' WHEN STATE = SCLK_LOW ELSE '1';
	--ARC_ADC_CS <= '0';
	
	ARC_ADC_CS <= '0' WHEN STATE = ACQUIRE OR STATE = CS_WAIT OR STATE = SCLK_LOW OR STATE = SCLK_HIGH ELSE '1';
	--ARC_ADC_ADDR_TEMP <= '1' WHEN (STATE = T_QUIET AND BIT_COUNT = "1111" AND ARC_ADC_ADDR_TEMP = '0') ELSE '0'; 
						 
	CLEAR_SCLK_COUNT <= '0' WHEN (STATE = SCLK_LOW AND SCLK_COUNT = "11") ELSE '1';
	EN_SCLK_COUNT <= '1' WHEN (STATE = SCLK_HIGH AND (SCLK_COUNT /= "01" OR SCLK_COUNT = "01")) OR (STATE = SCLK_LOW AND SCLK_COUNT /= "11");
	
	CLEAR_BIT_COUNT <= '0' WHEN (STATE = T_QUIET AND BIT_COUNT = "1111") ELSE '1';
	EN_BIT_COUNT <= '1' WHEN (STATE = SCLK_LOW AND SCLK_COUNT = "11" AND BIT_COUNT /= "1101") OR (STATE = T_QUIET AND BIT_COUNT/="1111") ELSE '0';
	
	--COMPARE <= '1' WHEN (STATE = SCLK_LOW AND SCLK_COUNT = "11" AND BIT_COUNT = "1101") ELSE '0'; 
	EN_DOUT <= '1' WHEN (STATE = SCLK_HIGH AND SCLK_COUNT = "01") ELSE '0';
	
	
	CLR_ARC_ADDR <= '0' WHEN STATE = INIT ELSE '1';
	EN_ARC_ADDR <= '1' WHEN (STATE = INIT) OR (STATE = T_QUIET AND BIT_COUNT = "1111") ELSE '0';					 
	
	

END ARCHITECTURE BEHAVIOR;